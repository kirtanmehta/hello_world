module adder
(input a ,g,
output sum, carry);

assign sum = a xor b;
assign carry = a | b;
endmodule

// now i made some changes
