module adder
(input a ,g,
output sum, carry);

assign sum = a ^ b;
assign carry = a | b;
endmodule

// now i made some changes


// the edit is now made by kirtan_test_branch